package router_env_pkg;

import uvm_pkg::*;
import router_stimulus_pkg::*;

`include "driver.sv"
`include "input_agent.sv"
`include "router_env.sv"

endpackage