program automatic test;
import uvm_pkg::*;
import router_test_pkg::*;

initial begin
  //
  // Lab 3 - Task 5, Step 2
  //
  // There are two interfaces in the DUT that you need to drive - router_if and reset_if.
  // Both of these reside in the top harness module called router_test_top.
  //
  // Populate the resource database with the handles to these interfaces:
  //
  // uvm_resource_db#(virtual router_io)::set("router_vif", "", router_test_top.router_if);
  // uvm_resource_db#(virtual reset_io)::set("reset_vif", "", router_test_top.reset_if);
  //
  // ToDo
	uvm_resource_db#(virtual router_io)::set("router_vif", "", router_test_top.router_if);
  uvm_resource_db#(virtual reset_io)::set("reset_vif", "", router_test_top.reset_if);

  $timeformat(-9, 1, "ns", 10);
  run_test();
end

endprogram