bind fifo fifo_sva 
i_fifo_bind
  (.*);
